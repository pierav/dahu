/* Config file */

package C;
    parameter int XLEN = 64;
endpackage
